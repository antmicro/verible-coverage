// Include whitespace around keywords and binary operators

parameter int I=1+2;
