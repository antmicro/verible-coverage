// begin must be on the same line as the preceding keyword and end the line

module begin_newline;
always_ff @(posedge clk)
begin end
endmodule
