// Each file should have only one module

module one_file_per_module;
// module name must be the same as file name
endmodule
module second;
endmodule
