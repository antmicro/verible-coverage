// For multiple items on a line, one space must separate the comma and the
// next character
module space_after_comma;
  int a,b,c;
endmodule
