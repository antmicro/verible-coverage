// Include whitespace around keywords and binary operators

module whitespace_keywords;endmodule
