// Line wraps should indent by four spaces
// This is the line length test after formatter

// verilog_syntax: parse-as-module-body
assign x = f;
assign lllllllllllllllllll[1111111111
  ] = aaaaaaaaaaa[4444444].ffffffffffffff.gggggggggggg.hhhhhhhhhhh.wwwww[555555].zzzzzzzzzz;
