// end must start a new line

module end_newline;
always @(posedge clk) begin
end endmodule
