// Style guide mandates two spaces per indent for all paired keywords.
class foo;
    function int validate();
    endfunction
endclass
